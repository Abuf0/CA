module efuse_rw_ctrl#(
    parameter NW = 64,
    parameter NR = 64
)(

);
endmodule