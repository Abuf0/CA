module efuse_write#(
    parameter NW = 64
)(

);
endmodule